
-- Modificado por Luis Jacobo �lvarez Ruiz de Ojeda el 7/7/2005 para evitar los errores que se
-- produc�an al intentar la simulaci�n funcional (y la temporal en ocasiones), debidos a la
-- definici�n del paquete "constants"

-- Modificado por Luis Jacobo �lvarez Ruiz de Ojeda el 17/10/2005 para evitar los avisos ("warnings" que se
-- produc�an al realizar la sintesis en Foundation ISE 7.1

library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package	constants is
	type TPicoType is ( pbtI, pbtII, pbt3, pbtS ) ;
	constant PicoType : TPicoType := pbt3 ;
	function ADDRSIZE return natural ;
	function INSTSIZE return natural ;
	function JADDRSIZE return natural ;
	function JDATASIZE return natural ;
end package ;

package body constants is
	function ADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 10 ;
		when pbt3 => return 10 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function INSTSIZE return natural is 
	begin
		case PicoType is
		when pbtI => return 16 ;
		when pbtII => return 18 ;
		when pbt3 => return 18 ;
		when pbtS => return 18 ;
		end case ;
	end ;
	function JADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 9 ;
		when pbtII => return 11 ;
		when pbt3 => return 11 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function JDATASIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 9 ;
		when pbt3 => return 9 ;
		when pbtS => return 20 ;
		end case ;
	end ;
end package body ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

-- La primera modificaci�n es poner la declaraci�n del uso del paquete "constants" antes de la de
-- la biblioteca "unisim", e indicar expresamente que el paquete pertenece a la biblioteca "work"
-- Este cambio es el que soluciona los problemas que se produc�an al intentar hacer
-- la simulaci�n temporal ("Post Map" y "Post Place & Route")
library work;
use work.constants.all;

library unisim ;
use unisim.vcomponents.all ;

entity picocode is
    port ( 
        clk : in std_logic ;
-- La segunda modificaci�n es eliminar la declaraci�n de la se�al de salida "reset", que en realidad no se utiliza
-- en este fichero sino en el correspondiente a la memoria de programa que se puede modificar via "Boundary Scan"	 
--        reset : out std_logic ;
        address : in std_logic_vector( ADDRSIZE - 1 downto 0 ) ;
        instruction : out std_logic_vector( INSTSIZE - 1 downto 0 )
    ) ;
end entity picocode ;

architecture mix of picocode is
    
-- La tercera modificaci�n es eliminar la declaraci�n del componente "jtag_shifter" que no se usa en
-- este fichero sino en el correspondiente a la memoria de programa que se puede modificar via "Boundary Scan"	 
--	 component jtag_shifter is
--        port ( 
--			clk : in std_logic ;
--			user1 : out std_logic ;
--            write : out std_logic ;
--            addr : out std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
--            data : out std_logic_vector( JDATASIZE - 1 downto 0 )
--        ) ;
--    end component ;

    signal jaddr : std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
    signal jdata : std_logic_vector( JDATASIZE - 1 downto 0 ) ;
    signal juser1 : std_logic ;
    signal jwrite : std_logic ;

-- La cuarta modificacion (del 17/10/2005) es eliminar la declaracion y asignacion de valores a todos los atributos
-- de inicializacion de las memorias BRAM, pues en Foundation ISE 7.1 se inicializan mediante el uso de "generic"
-- Ya no he dejado dichas l�neas en este fichero

begin

-- La quinta modificaci�n es sustituir en toda la descripci�n de la arquitectura las llamadas
-- a las funciones del paquete "constants" por los valores concretos que deben tomar en cada caso
-- Este cambio es el que soluciona los errores qe se produc�an al intentar hacer la simulaci�n funcional ("Behavioral")

	I18 : if (PicoType = pbtII) or (PicoType = pbt3) generate
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
					-- Modificaci�n del 8/3/2007
					-- Aqui hubo que a�adir estos par�metros para que no diese warnings en la versi�n ISE 8.2
					INIT_A => ('0' & X"00"), --  Value of output RAM registers on Port A at startup
					INIT_B => ("00" & X"0000"), --  Value of output RAM registers on Port B at startup
					SRVAL_A => ('0' & X"00"), --  Port A ouput value upon SSR assertion
					SRVAL_B => ("00" & X"0000"), --  Port B ouput value upon SSR assertion
					WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
					WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
					SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 			  
					-- Fin de la modificaci�n del 8/3/2007
	            INIT_00 => X"4803030002000500400BC001CA005006480148030B010A000901073D0656042E",
	            INIT_01 => X"48014803823085305C334002D010410140025819510041024001CB01500F4801",
	            INIT_02 => X"48014803C402502A48014803C202502648014803C702502248014803C602501E",
	            INIT_03 => X"000000000000403705008201401C5C334002503A450A8501C0028001C502502E",
	            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3F => X"400C000000000000000000000000000000000000000000000000000000000000",
	            INITP_00 => X"00000000000000000000000000000000031F757B4B4B4B4B45D4342D00FB4000",
	            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000"
	        )
	        port map (
	            DIB => "0000000000000000",
	            DIPB => "00",
	            ENB => '1',
	            WEB => '0',
	            SSRB => '0',
	            CLKB => clk,
	            ADDRB => address,
	            DOB => instruction( 18 - 3 downto 0 ),		-- Aqu� se sustituy� la funci�n por su valor concreto
	            DOPB => instruction( 18 - 1 downto 18 - 2 ),		-- Aqu� se sustituy� la funci�n por su valor concreto
	            DIA => jdata( 9 - 2 downto 0 ),		-- Aqu� se sustituy� la funci�n por su valor concreto
	            DIPA => jdata( 9 - 1 downto 9 - 1 ),		-- Aqu� se sustituy� la funci�n por su valor concreto
	            ENA => juser1,
	            WEA => jwrite,
	            SSRA => '0',
	            CLKA => clk,
	            ADDRA => jaddr,
	            DOA => open,
	            DOPA => open 
	        ) ;
	end generate ;

	I16 : if PicoType = pbtI generate
	begin
	    bram : component RAMB4_S8_S16
	        generic map (
	            INIT_00 => X"4803030002000500400BC001CA005006480148030B010A000901073D0656042E",
	            INIT_01 => X"48014803823085305C334002D010410140025819510041024001CB01500F4801",
	            INIT_02 => X"48014803C402502A48014803C202502648014803C702502248014803C602501E",
	            INIT_03 => X"000000000000403705008201401C5C334002503A450A8501C0028001C502502E",
	            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIB => "0000000000000000",  
				ENB => '1', 
				WEB => '0',
				RSTB =>	'0',
				CLKB => clk,
				ADDRB => address,
				DOB => instruction( 16 - 1 downto 0 ),  		-- Aqu� se sustituy� la funci�n por su valor concreto
				DIA => jdata( 8 - 1 downto 0 ),   		-- Aqu� se sustituy� la funci�n por su valor concreto
				ENA => juser1, 
				WEA => jwrite,
				RSTA => '0',
				CLKA => clk,
				ADDRA => jaddr,
				DOA => open  
			) ; 
	end generate ;

	I20 : if PicoType = pbtS generate
		signal data_out : std_logic_vector( 3 downto 0 ) ;
	begin
	    ram_1 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0003013313111323102310231023102310113110031002310000332310000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"3000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => data_out,  
				DIB => jdata( 20 - 1 downto 16 ),   		-- Aqu� se sustituy� la funci�n por su valor concreto
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
			-- loose top 2 bits
			instruction( 17 downto 16 ) <= data_out( 1 downto 0 ) ;

	    ram_2 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"000408454548C8C544C544C544C544C5448854D445544C5440004CC544000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"4000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 15 downto 12 ),  
				DIB => jdata( 15 downto 12 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_3 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0000520C0055005088408820887088608825C00108110B08832500A088BA9764",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 11 downto 8 ),  
				DIB => jdata( 11 downto 8 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_4 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0003001303000002000200020002000100333010010000000000000000000352",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 7 downto 4 ),  
				DIB => jdata( 7 downto 4 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_5 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"000701C32AA1212E132A13261322132E13003201290211F13000B10613101D6E",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"C000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 3 downto 0 ),  
				DIB => jdata( 3 downto 0 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
	end generate ;

	jdata <= ( others => '0' ) ;
	jaddr <= ( others => '0' ) ;
	juser1 <= '0' ;
	jwrite <= '0' ;
end architecture mix ;
